module reg(dataIn,reset,En,dataOut);



endmodule